ENTITY MAC_SNACKS IS
    PORT(CLK, INSERTING, SELECT_I, CANCEL: IN BIT;
        VALUE: IN BIT_VECTOR(3 DOWNTO 0);
        COD_PROD: IN BIT_VECTOR(1 DOWNTO 0);
        IS_RELEASE: OUT BIT;
        REMAINING_MONEY: OUT BIT_VECTOR(3 DOWNTO 0));
END MAC_SNACKS;

ARCHITECTURE LOGIC OF MAC_SNACKS IS

COMPONENT CON_BLOCK IS
    PORT(CLK, INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL: IN BIT;
        IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM: OUT BIT);
END COMPONENT;

COMPONENT OP_BLOCK IS
    PORT (VALUE: IN BIT_VECTOR(3 DOWNTO 0);
        COD_PROD: IN BIT_VECTOR(1 DOWNTO 0);
        ACC_LD, ACC_CLR, S_RM, RM_LD, RM_CLR, CLK: IN BIT;
        REMAINING_MONEY: OUT BIT_VECTOR(3 DOWNTO 0);
        GTEQ_VALUE, LT_16: OUT BIT
    );
END COMPONENT;

SIGNAL ACC_LD, ACC_CLR, RM_LD, RM_CLR, S_RM, GTEQ_VALUE, LT_16: BIT;

BEGIN 

    BLOCO_DE_CONTROLE: CON_BLOCK PORT MAP(CLK, INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL, IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM);
    BLOCO_OPERACIONAL: OP_BLOCK PORT MAP(VALUE, COD_PROD, ACC_LD, ACC_CLR, S_RM, RM_LD, RM_CLR, CLK, REMAINING_MONEY, GTEQ_VALUE, LT_16);

END LOGIC;