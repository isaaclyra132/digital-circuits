library ieee ;
use ieee.std_logic_1164.all;

ENTITY MDE_B IS
    PORT(CLK, RST, INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL: IN STD_LOGIC;
        IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM: OUT STD_LOGIC);
END MDE_B;

ARCHITECTURE LOGIC OF MDE_B IS
    TYPE STATE_TYPE is (INICIO, ESPERA, SOMA, ESCOLHE, LIBERA, CANCELA);
    SIGNAL Y_PRESENT, Y_NEXT: STATE_TYPE;
BEGIN
    PROCESS(INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL, Y_PRESENT)
    BEGIN
        CASE Y_PRESENT IS
        WHEN INICIO =>
            Y_NEXT <= ESPERA;
        WHEN ESPERA =>
            IF (INSERTING = '0' AND SELECT_I = '0' AND CANCEL = '0') THEN Y_NEXT <= ESPERA;
            ELSIF (INSERTING = '1' AND LT_16 = '1' AND CANCEL = '0') THEN Y_NEXT <= SOMA;
            ELSIF (INSERTING = '0' AND SELECT_I = '1' AND CANCEL = '0') THEN Y_NEXT <= ESCOLHE;
            ELSIF (CANCEL = '1') THEN Y_NEXT <= CANCELA;
            END IF;
        WHEN SOMA =>
            Y_NEXT <= ESPERA;
        WHEN ESCOLHE =>
            IF (GTEQ_VALUE = '0') THEN Y_NEXT <= ESPERA;
            ELSIF (GTEQ_VALUE = '1') THEN Y_NEXT <= LIBERA;
            END IF;
        WHEN LIBERA =>
            Y_NEXT <= INICIO;
        WHEN CANCELA =>
            Y_NEXT <= INICIO;
        END CASE;
    END PROCESS;

    PROCESS (CLK, RST)
    BEGIN
        IF RST = '1' THEN
            Y_PRESENT <= INICIO;
        ELSIF (CLK'event AND CLK = '1') THEN
            Y_PRESENT <= Y_NEXT;
        END IF;
    END PROCESS;

    IS_RELEASE <= '1' WHEN Y_PRESENT = LIBERA ELSE '0';
    ACC_CLR <= '1' WHEN Y_PRESENT = INICIO ELSE '0';
    ACC_LD <= '1' WHEN Y_PRESENT = SOMA ELSE '0';
    RM_CLR <= '1' WHEN Y_PRESENT = INICIO ELSE '0';
    RM_LD <= '1' WHEN (Y_PRESENT = LIBERA OR Y_PRESENT = CANCELA) ELSE '0';
    S_RM <= '1' WHEN Y_PRESENT = LIBERA ELSE '0';
    
END LOGIC;