ENTITY MDE IS
    PORT(Q2, Q1, Q0, INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL: IN BIT;
        D2, D1, D0, IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM: OUT BIT);
END MDE;

ARCHITECTURE LOGIC OF MDE IS

BEGIN

D2 <= (NOT Q2 AND NOT Q1 AND Q0 AND NOT INSERTING AND NOT SELECT_I AND NOT LT_16 AND NOT GTEQ_VALUE AND CANCEL)
    OR (NOT Q2 AND Q1 AND Q0 AND NOT INSERTING AND NOT SELECT_I AND NOT LT_16 AND GTEQ_VALUE AND NOT CANCEL);
D1 <= (NOT Q2 AND NOT Q1 AND Q0 AND NOT INSERTING AND SELECT_I AND NOT CANCEL)
    OR (NOT Q2 AND NOT Q1 AND Q0 AND INSERTING AND LT_16 AND NOT CANCEL);
D0 <= (NOT Q2 AND NOT INSERTING AND NOT SELECT_I AND NOT LT_16 AND NOT GTEQ_VALUE AND NOT CANCEL)
    OR (NOT Q2 AND NOT Q1 AND Q0 AND NOT INSERTING AND NOT SELECT_I AND NOT LT_16 AND NOT GTEQ_VALUE)
    OR (NOT Q2 AND NOT Q1 AND Q0 AND NOT INSERTING AND NOT LT_16 AND NOT GTEQ_VALUE AND NOT CANCEL);
IS_RELEASE <= Q2 AND NOT Q1 AND NOT Q0;
ACC_CLR <= NOT Q2 AND NOT Q1 AND NOT Q0;
ACC_LD <= NOT Q2 AND Q1 AND NOT Q0;
RM_CLR <= NOT Q2 AND NOT Q1 AND NOT Q0;
RM_LD <= (Q2 AND NOT Q1 AND NOT Q0) OR (Q2 AND NOT Q1 AND Q0);
S_RM <= Q2 AND NOT Q1 AND NOT Q0;

END LOGIC;