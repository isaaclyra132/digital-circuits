ENTITY CON_BLOCK IS
    PORT(CLK, INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL: IN BIT;
        IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM: OUT BIT);
END CON_BLOCK;

ARCHITECTURE LOGIC OF CON_BLOCK IS

COMPONENT MDE IS
    PORT(Q2, Q1, Q0, INSERTING, SELECT_I, LT_16, GTEQ_VALUE, CANCEL: IN BIT;
        D2, D1, D0, IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM: OUT BIT);
END COMPONENT;

COMPONENT ffd IS
	port ( clk ,D ,P , C : IN BIT ;
		q : OUT BIT );
END COMPONENT ;

COMPONENT BS IS
    PORT(CLK, T: IN BIT;
        PRESS: OUT BIT);
END COMPONENT;

SIGNAL Q2, Q1, Q0, D2, D1, D0, PRESS_INSERTING, PRESS_SELECT, PRESS_CANCEL: BIT;

BEGIN

-- BOTÕES SÍNCRONOS
BUTTON_INSERTING: BS PORT MAP(CLK, INSERTING, PRESS_INSERTING);
BUTTON_SELECT: BS PORT MAP(CLK, SELECT_I, PRESS_SELECT);
BUTTON_CANCEL: BS PORT MAP(CLK, CANCEL, PRESS_CANCEL);

-- LÓGICA COMBINACIONAL DO BLOCO DE CONTROLE
LOGIC: MDE PORT MAP(Q2, Q1, Q0, PRESS_INSERTING, PRESS_SELECT, LT_16, GTEQ_VALUE, PRESS_CANCEL, D2, D1, D0, IS_RELEASE, ACC_CLR, ACC_LD, RM_CLR, RM_LD, S_RM);

-- REGISTRADORES DE ESTADO
REG_STATE_BIT0: ffd PORT MAP(CLK, D0, '1', '1', Q0);
REG_STATE_BIT1: ffd PORT MAP(CLK, D1, '1', '1', Q1);
REG_STATE_BIT2: ffd PORT MAP(CLK, D2, '1', '1', Q2);

END LOGIC;