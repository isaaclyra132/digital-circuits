ENTITY OP_BLOCK IS
    PORT (VALUE: IN BIT_VECTOR(3 DOWNTO 0);
        COD_PROD: IN BIT_VECTOR(1 DOWNTO 0);
        ACC_LD, ACC_CLR, S_RM, RM_LD, RM_CLR, CLK: IN BIT;
        REMAINING_MONEY: OUT BIT_VECTOR(3 DOWNTO 0);
        GTEQ_VALUE, LT_16: OUT BIT
    );
END OP_BLOCK;

ARCHITECTURE LOGIC OF OP_BLOCK IS

COMPONENT REG4 is
	port(A: in bit_vector(3 downto 0);
		ld, clk, clr: in bit;
		S: out bit_vector(3 downto 0));
end COMPONENT;

COMPONENT MUX41_4B IS
    PORT(I0, I1, I2, I3: IN BIT_VECTOR(3 DOWNTO 0);
        S: IN BIT_VECTOR(1 DOWNTO 0);
        O: OUT BIT_VECTOR(3 DOWNTO 0));
END COMPONENT;

COMPONENT MUX21_4B is
    port(I0, I1: in bit_vector(3 downto 0);
        S: in bit;
        O: out bit_vector(3 downto 0)
        );
end COMPONENT;

COMPONENT COMP_4B IS
  PORT(
      A, B: IN bit_vector(3 downto 0);
      LT: OUT BIT;
      EQ: OUT BIT;
      GT: OUT BIT
  );
END COMPONENT;

COMPONENT ADDER_4B is
    port (
        A, B: in bit_vector(3 downto 0);
        O: out bit_vector(3 downto 0);
        cout: out bit
    );
end COMPONENT;

COMPONENT SUB_4B is
    port (
        A, B: in bit_vector(3 downto 0);
        O: out bit_vector(3 downto 0);
        cout: out bit
    );
end COMPONENT;

SIGNAL PROD_VALUE0, PROD_VALUE1, PROD_VALUE2, PROD_VALUE3, VALUE_PROD0, VALUE_PROD1, VALUE_PROD2, 
        VALUE_PROD3, REG_OUT, ADD_RES, SUB_RES, PRODUCT_VALUE, RM_MUX: BIT_VECTOR(3 DOWNTO 0);
SIGNAL COMP_OUT: BIT_VECTOR(1 DOWNTO 0);
SIGNAL LIXO: BIT_VECTOR(4 DOWNTO 0);

BEGIN

-- VALORES DOS PRODUTOS E REGISTRADORES
PROD_VALUE0 <= "0101";
PROD_VALUE1 <= "1010";
PROD_VALUE2 <= "1000";
PROD_VALUE3 <= "0101";
REG_PROD0: REG4 PORT MAP(PROD_VALUE0, '1', CLK, '1', VALUE_PROD0);
REG_PROD1: REG4 PORT MAP(PROD_VALUE1, '1', CLK, '1', VALUE_PROD1);
REG_PROD2: REG4 PORT MAP(PROD_VALUE2, '1', CLK, '1', VALUE_PROD2);
REG_PROD3: REG4 PORT MAP(PROD_VALUE3, '1', CLK, '1', VALUE_PROD3);

-- MUX SELETOR DO PRODUTO
MUX_PROD: MUX41_4B PORT MAP(VALUE_PROD0, VALUE_PROD1, VALUE_PROD2, VALUE_PROD3, COD_PROD, PRODUCT_VALUE);

-- SOMADOR E REGISTRADOR
SOMA: ADDER_4B PORT MAP(VALUE, REG_OUT, ADD_RES, LIXO(0));
REG_ACC: REG4 PORT MAP(ADD_RES, ACC_LD, CLK, ACC_CLR, REG_OUT);

-- COMPARADOR DO ACUMULADOR X VALOR DO PRODUTO SELECIONADO
COMP_MONEY: COMP_4B PORT MAP(REG_OUT, PRODUCT_VALUE, LIXO(1), COMP_OUT(0), COMP_OUT(1));
GTEQ_VALUE <= COMP_OUT(0) OR COMP_OUT(1);

-- SUBTRAÇÃO
SUB_REM: SUB_4B PORT MAP(REG_OUT, PRODUCT_VALUE, SUB_RES, LIXO(2));

-- MUX SELETOR DO REMAINING MONEY
MUX_REM: MUX21_4B PORT MAP(REG_OUT, SUB_RES, S_RM, RM_MUX);

-- REGISTRADOR DE REMAINING MONEY
RESTO: REG4 PORT MAP(RM_MUX, RM_LD, CLK, RM_CLR, REMAINING_MONEY);

-- DEFINIÇÃO DE LT_16
COMP_LT: COMP_4B PORT MAP(ADD_RES, "1111", LT_16, LIXO(3), LIXO(4));

END LOGIC;